`timescale 1ns / 1ps
module CU (
    input wire[5:0] opcode,
    output wire[8:0] cu_out
);
    
endmodule